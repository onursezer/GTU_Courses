library verilog;
use verilog.vl_types.all;
entity sezer_onur_121044074 is
    port(
        result          : out    vl_logic_vector(31 downto 0)
    );
end sezer_onur_121044074;
