library verilog;
use verilog.vl_types.all;
entity main is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end main;
