library verilog;
use verilog.vl_types.all;
entity test_main is
end test_main;
